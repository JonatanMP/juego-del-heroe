module contador (
    
);

endmodule //contador